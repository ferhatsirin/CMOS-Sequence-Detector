magic
tech scmos
timestamp 1578742312
<< nwell >>
rect -221 247 -188 276
rect -162 251 -105 278
rect -70 247 -37 276
rect -11 239 31 266
rect 70 247 103 276
rect -224 181 -184 209
rect -166 153 -133 182
rect -73 181 -33 209
rect -13 181 18 182
rect 67 181 107 209
rect -15 153 18 181
rect 125 153 158 182
rect -221 105 -181 134
rect -168 87 -128 115
rect -70 105 -30 134
rect -17 87 23 115
rect 70 105 110 134
rect 123 87 163 115
rect -223 36 -183 64
rect -168 18 -128 45
rect -72 36 -32 64
rect -8 12 16 39
rect 68 36 108 64
<< ntransistor >>
rect -210 224 -208 229
rect -202 224 -200 229
rect -59 224 -57 229
rect -51 224 -49 229
rect -151 212 -149 217
rect -143 212 -141 217
rect -135 212 -133 217
rect -127 212 -125 217
rect -119 212 -117 217
rect 81 224 83 229
rect 89 224 91 229
rect 1 201 3 206
rect 9 201 11 206
rect 17 201 19 206
rect -213 153 -211 158
rect -205 153 -203 158
rect -197 153 -195 158
rect -62 153 -60 158
rect -54 153 -52 158
rect -46 153 -44 158
rect 78 153 80 158
rect 86 153 88 158
rect 94 153 96 158
rect -155 130 -153 135
rect -147 130 -145 135
rect -4 130 -2 135
rect 4 130 6 135
rect 136 130 138 135
rect 144 130 146 135
rect -210 79 -208 84
rect -202 79 -200 84
rect -194 79 -192 84
rect -59 79 -57 84
rect -51 79 -49 84
rect -43 79 -41 84
rect 81 79 83 84
rect 89 79 91 84
rect 97 79 99 84
rect -157 59 -155 64
rect -149 59 -147 64
rect -141 59 -139 64
rect -6 59 -4 64
rect 2 59 4 64
rect 10 59 12 64
rect 134 59 136 64
rect 142 59 144 64
rect 150 59 152 64
rect -212 8 -210 13
rect -204 8 -202 13
rect -196 8 -194 13
rect -61 8 -59 13
rect -53 8 -51 13
rect -45 8 -43 13
rect -157 2 -155 7
rect -149 2 -147 7
rect -141 2 -139 7
rect 79 8 81 13
rect 87 8 89 13
rect 95 8 97 13
rect 3 1 5 6
<< ptransistor >>
rect -210 253 -208 263
rect -202 253 -200 263
rect -151 257 -149 267
rect -143 257 -141 267
rect -135 257 -133 267
rect -127 257 -125 267
rect -119 257 -117 267
rect -59 253 -57 263
rect -51 253 -49 263
rect 1 245 3 255
rect 9 245 11 255
rect 17 245 19 255
rect 81 253 83 263
rect 89 253 91 263
rect -213 188 -211 198
rect -205 188 -203 198
rect -197 188 -195 198
rect -62 188 -60 198
rect -54 188 -52 198
rect -46 188 -44 198
rect 78 188 80 198
rect 86 188 88 198
rect 94 188 96 198
rect -155 159 -153 169
rect -147 159 -145 169
rect -4 159 -2 169
rect 4 159 6 169
rect 136 159 138 169
rect 144 159 146 169
rect -210 111 -208 121
rect -202 111 -200 121
rect -194 111 -192 121
rect -59 111 -57 121
rect -51 111 -49 121
rect -43 111 -41 121
rect -157 94 -155 104
rect -149 94 -147 104
rect -141 94 -139 104
rect 81 111 83 121
rect 89 111 91 121
rect 97 111 99 121
rect -6 94 -4 104
rect 2 94 4 104
rect 10 94 12 104
rect 134 94 136 104
rect 142 94 144 104
rect 150 94 152 104
rect -212 43 -210 53
rect -204 43 -202 53
rect -196 43 -194 53
rect -61 43 -59 53
rect -53 43 -51 53
rect -45 43 -43 53
rect -157 24 -155 34
rect -149 24 -147 34
rect -141 24 -139 34
rect 79 43 81 53
rect 87 43 89 53
rect 95 43 97 53
rect 3 18 5 28
<< ndiffusion >>
rect -211 224 -210 229
rect -208 224 -202 229
rect -200 224 -199 229
rect -60 224 -59 229
rect -57 224 -51 229
rect -49 224 -48 229
rect -152 212 -151 217
rect -149 212 -148 217
rect -144 212 -143 217
rect -141 212 -140 217
rect -136 212 -135 217
rect -133 212 -132 217
rect -128 212 -127 217
rect -125 212 -124 217
rect -120 212 -119 217
rect -117 212 -116 217
rect 80 224 81 229
rect 83 224 89 229
rect 91 224 92 229
rect 0 201 1 206
rect 3 201 9 206
rect 11 201 12 206
rect 16 201 17 206
rect 19 201 20 206
rect -214 153 -213 158
rect -211 153 -205 158
rect -203 153 -197 158
rect -195 153 -194 158
rect -63 153 -62 158
rect -60 153 -54 158
rect -52 153 -46 158
rect -44 153 -43 158
rect 77 153 78 158
rect 80 153 86 158
rect 88 153 94 158
rect 96 153 97 158
rect -156 130 -155 135
rect -153 130 -147 135
rect -145 130 -144 135
rect -5 130 -4 135
rect -2 130 4 135
rect 6 130 7 135
rect 135 130 136 135
rect 138 130 144 135
rect 146 130 147 135
rect -211 79 -210 84
rect -208 79 -202 84
rect -200 79 -194 84
rect -192 79 -191 84
rect -60 79 -59 84
rect -57 79 -51 84
rect -49 79 -43 84
rect -41 79 -40 84
rect 80 79 81 84
rect 83 79 89 84
rect 91 79 97 84
rect 99 79 100 84
rect -158 59 -157 64
rect -155 59 -149 64
rect -147 59 -141 64
rect -139 59 -138 64
rect -7 59 -6 64
rect -4 59 2 64
rect 4 59 10 64
rect 12 59 13 64
rect 133 59 134 64
rect 136 59 142 64
rect 144 59 150 64
rect 152 59 153 64
rect -213 8 -212 13
rect -210 8 -204 13
rect -202 8 -196 13
rect -194 8 -193 13
rect -62 8 -61 13
rect -59 8 -53 13
rect -51 8 -45 13
rect -43 8 -42 13
rect -158 2 -157 7
rect -155 2 -154 7
rect -150 2 -149 7
rect -147 2 -146 7
rect -142 2 -141 7
rect -139 2 -138 7
rect 78 8 79 13
rect 81 8 87 13
rect 89 8 95 13
rect 97 8 98 13
rect 2 1 3 6
rect 5 1 6 6
<< pdiffusion >>
rect -211 253 -210 263
rect -208 253 -207 263
rect -203 253 -202 263
rect -200 253 -199 263
rect -152 257 -151 267
rect -149 257 -143 267
rect -141 257 -135 267
rect -133 257 -132 267
rect -128 257 -127 267
rect -125 257 -119 267
rect -117 257 -116 267
rect -60 253 -59 263
rect -57 253 -56 263
rect -52 253 -51 263
rect -49 253 -48 263
rect 0 245 1 255
rect 3 245 4 255
rect 8 245 9 255
rect 11 245 12 255
rect 16 245 17 255
rect 19 245 20 255
rect 80 253 81 263
rect 83 253 84 263
rect 88 253 89 263
rect 91 253 92 263
rect -214 188 -213 198
rect -211 188 -210 198
rect -206 188 -205 198
rect -203 188 -202 198
rect -198 188 -197 198
rect -195 188 -194 198
rect -63 188 -62 198
rect -60 188 -59 198
rect -55 188 -54 198
rect -52 188 -51 198
rect -47 188 -46 198
rect -44 188 -43 198
rect 77 188 78 198
rect 80 188 81 198
rect 85 188 86 198
rect 88 188 89 198
rect 93 188 94 198
rect 96 188 97 198
rect -156 159 -155 169
rect -153 159 -152 169
rect -148 159 -147 169
rect -145 159 -144 169
rect -5 159 -4 169
rect -2 159 -1 169
rect 3 159 4 169
rect 6 159 7 169
rect 135 159 136 169
rect 138 159 139 169
rect 143 159 144 169
rect 146 159 147 169
rect -211 111 -210 121
rect -208 111 -207 121
rect -203 111 -202 121
rect -200 111 -199 121
rect -195 111 -194 121
rect -192 111 -191 121
rect -60 111 -59 121
rect -57 111 -56 121
rect -52 111 -51 121
rect -49 111 -48 121
rect -44 111 -43 121
rect -41 111 -40 121
rect -158 94 -157 104
rect -155 94 -154 104
rect -150 94 -149 104
rect -147 94 -146 104
rect -142 94 -141 104
rect -139 94 -138 104
rect 80 111 81 121
rect 83 111 84 121
rect 88 111 89 121
rect 91 111 92 121
rect 96 111 97 121
rect 99 111 100 121
rect -7 94 -6 104
rect -4 94 -3 104
rect 1 94 2 104
rect 4 94 5 104
rect 9 94 10 104
rect 12 94 13 104
rect 133 94 134 104
rect 136 94 137 104
rect 141 94 142 104
rect 144 94 145 104
rect 149 94 150 104
rect 152 94 153 104
rect -213 43 -212 53
rect -210 43 -209 53
rect -205 43 -204 53
rect -202 43 -201 53
rect -197 43 -196 53
rect -194 43 -193 53
rect -62 43 -61 53
rect -59 43 -58 53
rect -54 43 -53 53
rect -51 43 -50 53
rect -46 43 -45 53
rect -43 43 -42 53
rect -158 24 -157 34
rect -155 24 -149 34
rect -147 24 -141 34
rect -139 24 -138 34
rect 78 43 79 53
rect 81 43 82 53
rect 86 43 87 53
rect 89 43 90 53
rect 94 43 95 53
rect 97 43 98 53
rect 2 18 3 28
rect 5 18 6 28
<< ndcontact >>
rect -215 224 -211 229
rect -199 224 -194 229
rect -64 224 -60 229
rect -48 224 -43 229
rect -156 212 -152 217
rect -148 212 -144 217
rect -140 212 -136 217
rect -132 212 -128 217
rect -124 212 -120 217
rect -116 212 -112 217
rect 76 224 80 229
rect 92 224 97 229
rect -4 201 0 206
rect 12 201 16 206
rect 20 201 24 206
rect -218 153 -214 158
rect -194 153 -189 158
rect -67 153 -63 158
rect -43 153 -38 158
rect 73 153 77 158
rect 97 153 102 158
rect -160 130 -156 135
rect -144 130 -139 135
rect -9 130 -5 135
rect 7 130 12 135
rect 131 130 135 135
rect 147 130 152 135
rect -215 79 -211 84
rect -191 79 -186 84
rect -64 79 -60 84
rect -40 79 -35 84
rect 76 79 80 84
rect 100 79 105 84
rect -162 59 -158 64
rect -138 59 -133 64
rect -11 59 -7 64
rect 13 59 18 64
rect 129 59 133 64
rect 153 59 158 64
rect -217 8 -213 13
rect -193 8 -188 13
rect -66 8 -62 13
rect -42 8 -37 13
rect -162 2 -158 7
rect -154 2 -150 7
rect -146 2 -142 7
rect -138 2 -134 7
rect 74 8 78 13
rect 98 8 103 13
rect -2 1 2 6
rect 6 1 10 6
<< pdcontact >>
rect -215 253 -211 263
rect -207 253 -203 263
rect -199 253 -195 263
rect -156 257 -152 267
rect -132 257 -128 267
rect -116 257 -112 267
rect -64 253 -60 263
rect -56 253 -52 263
rect -48 253 -44 263
rect -4 245 0 255
rect 4 245 8 255
rect 12 245 16 255
rect 20 245 24 255
rect 76 253 80 263
rect 84 253 88 263
rect 92 253 96 263
rect -218 188 -214 198
rect -210 188 -206 198
rect -202 188 -198 198
rect -194 188 -190 198
rect -67 188 -63 198
rect -59 188 -55 198
rect -51 188 -47 198
rect -43 188 -39 198
rect 73 188 77 198
rect 81 188 85 198
rect 89 188 93 198
rect 97 188 101 198
rect -160 159 -156 169
rect -152 159 -148 169
rect -144 159 -140 169
rect -9 159 -5 169
rect -1 159 3 169
rect 7 159 11 169
rect 131 159 135 169
rect 139 159 143 169
rect 147 159 151 169
rect -215 111 -211 121
rect -207 111 -203 121
rect -199 111 -195 121
rect -191 111 -187 121
rect -64 111 -60 121
rect -56 111 -52 121
rect -48 111 -44 121
rect -40 111 -36 121
rect -162 94 -158 104
rect -154 94 -150 104
rect -146 94 -142 104
rect -138 94 -134 104
rect 76 111 80 121
rect 84 111 88 121
rect 92 111 96 121
rect 100 111 104 121
rect -11 94 -7 104
rect -3 94 1 104
rect 5 94 9 104
rect 13 94 17 104
rect 129 94 133 104
rect 137 94 141 104
rect 145 94 149 104
rect 153 94 157 104
rect -217 43 -213 53
rect -209 43 -205 53
rect -201 43 -197 53
rect -193 43 -189 53
rect -66 43 -62 53
rect -58 43 -54 53
rect -50 43 -46 53
rect -42 43 -38 53
rect -162 24 -158 34
rect -138 24 -134 34
rect 74 43 78 53
rect 82 43 86 53
rect 90 43 94 53
rect 98 43 102 53
rect -2 18 2 28
rect 6 18 10 28
<< psubstratepcontact >>
rect -215 215 -211 219
rect -207 215 -203 219
rect -199 215 -195 219
rect -64 215 -60 219
rect -56 215 -52 219
rect -48 215 -44 219
rect 76 215 80 219
rect 84 215 88 219
rect 92 215 96 219
rect -4 193 0 197
rect 4 193 8 197
rect 12 193 16 197
rect 20 193 24 197
rect -218 145 -214 149
rect -210 145 -206 149
rect -202 145 -198 149
rect -194 145 -190 149
rect -67 145 -63 149
rect -59 145 -55 149
rect -51 145 -47 149
rect -43 145 -39 149
rect 73 145 77 149
rect 81 145 85 149
rect 89 145 93 149
rect 97 145 101 149
rect -160 121 -156 125
rect -152 121 -148 125
rect -144 121 -140 125
rect -9 121 -5 125
rect -1 121 3 125
rect 7 121 11 125
rect 131 121 135 125
rect 139 121 143 125
rect 147 121 151 125
rect -215 70 -211 74
rect -207 70 -203 74
rect -199 70 -195 74
rect -191 70 -187 74
rect -64 70 -60 74
rect -56 70 -52 74
rect -48 70 -44 74
rect -40 70 -36 74
rect 76 70 80 74
rect 84 70 88 74
rect 92 70 96 74
rect 100 70 104 74
rect -162 51 -158 55
rect -154 51 -150 55
rect -146 51 -142 55
rect -138 51 -134 55
rect -11 51 -7 55
rect -3 51 1 55
rect 5 51 9 55
rect 13 51 17 55
rect 129 51 133 55
rect 137 51 141 55
rect 145 51 149 55
rect 153 51 157 55
rect -217 0 -213 4
rect -209 0 -205 4
rect -201 0 -197 4
rect -193 0 -189 4
rect -162 -6 -158 -2
rect -154 -6 -150 -2
rect -66 0 -62 4
rect -58 0 -54 4
rect -50 0 -46 4
rect -42 0 -38 4
rect 74 0 78 4
rect 82 0 86 4
rect 90 0 94 4
rect 98 0 102 4
rect -146 -6 -142 -2
rect -138 -6 -134 -2
rect -2 -7 2 -3
rect 6 -7 10 -3
<< nsubstratencontact >>
rect -215 268 -211 272
rect -207 268 -203 272
rect -199 268 -195 272
rect -156 271 -152 275
rect -148 271 -144 275
rect -140 271 -136 275
rect -132 271 -128 275
rect -124 271 -120 275
rect -116 271 -112 275
rect -64 268 -60 272
rect -56 268 -52 272
rect -48 268 -44 272
rect -4 259 0 263
rect 4 259 8 263
rect 12 259 16 263
rect 20 259 24 263
rect 76 268 80 272
rect 84 268 88 272
rect 92 268 96 272
rect -218 202 -214 206
rect -210 202 -206 206
rect -202 202 -198 206
rect -194 202 -190 206
rect -156 199 -152 203
rect -148 199 -144 203
rect -140 199 -136 203
rect -132 199 -128 203
rect -124 199 -120 203
rect -116 199 -112 203
rect -67 202 -63 206
rect -59 202 -55 206
rect -51 202 -47 206
rect -43 202 -39 206
rect 73 202 77 206
rect 81 202 85 206
rect 89 202 93 206
rect 97 202 101 206
rect -160 174 -156 178
rect -152 174 -148 178
rect -144 174 -140 178
rect -9 174 -5 178
rect -1 174 3 178
rect 7 174 11 178
rect 131 174 135 178
rect 139 174 143 178
rect 147 174 151 178
rect -215 126 -211 130
rect -207 126 -203 130
rect -199 126 -195 130
rect -191 126 -187 130
rect -64 126 -60 130
rect -56 126 -52 130
rect -48 126 -44 130
rect -40 126 -36 130
rect 76 126 80 130
rect 84 126 88 130
rect 92 126 96 130
rect 100 126 104 130
rect -162 108 -158 112
rect -154 108 -150 112
rect -146 108 -142 112
rect -138 108 -134 112
rect -11 108 -7 112
rect -3 108 1 112
rect 5 108 9 112
rect 13 108 17 112
rect 129 108 133 112
rect 137 108 141 112
rect 145 108 149 112
rect 153 108 157 112
rect -217 57 -213 61
rect -209 57 -205 61
rect -201 57 -197 61
rect -193 57 -189 61
rect -66 57 -62 61
rect -58 57 -54 61
rect -50 57 -46 61
rect -42 57 -38 61
rect 74 57 78 61
rect 82 57 86 61
rect 90 57 94 61
rect 98 57 102 61
rect -162 38 -158 42
rect -154 38 -150 42
rect -146 38 -142 42
rect -138 38 -134 42
rect -2 32 2 36
rect 6 32 10 36
<< polysilicon >>
rect -151 267 -149 270
rect -143 267 -141 270
rect -135 267 -133 270
rect -127 267 -125 270
rect -119 267 -117 284
rect -95 272 -93 297
rect -210 263 -208 266
rect -202 263 -200 266
rect -231 237 -229 247
rect -210 244 -208 253
rect -210 229 -208 240
rect -202 237 -200 253
rect -202 229 -200 233
rect -151 231 -149 257
rect -143 252 -141 257
rect -210 221 -208 224
rect -202 221 -200 224
rect -151 217 -149 227
rect -143 217 -141 248
rect -135 245 -133 257
rect -135 217 -133 241
rect -127 238 -125 257
rect -127 217 -125 234
rect -119 217 -117 257
rect -81 237 -79 287
rect 45 272 47 293
rect -59 263 -57 266
rect -51 263 -49 266
rect 1 255 3 258
rect 9 255 11 258
rect 17 255 19 258
rect -59 244 -57 253
rect -59 229 -57 240
rect -51 237 -49 253
rect 1 234 3 245
rect -51 229 -49 233
rect -59 221 -57 224
rect -51 221 -49 224
rect -151 209 -149 212
rect -143 209 -141 212
rect -135 209 -133 212
rect -127 209 -125 212
rect -119 209 -117 212
rect 1 206 3 230
rect 9 227 11 245
rect 9 206 11 223
rect 17 220 19 245
rect 60 237 62 287
rect 81 263 83 266
rect 89 263 91 266
rect 81 244 83 253
rect 81 229 83 240
rect 89 237 91 253
rect 89 229 91 233
rect 81 221 83 224
rect 89 221 91 224
rect 17 206 19 216
rect -213 198 -211 201
rect -205 198 -203 201
rect -197 198 -195 201
rect -62 198 -60 201
rect -54 198 -52 201
rect -46 198 -44 201
rect 1 198 3 201
rect 9 198 11 201
rect 17 198 19 201
rect 78 198 80 201
rect 86 198 88 201
rect 94 198 96 201
rect -213 170 -211 188
rect -205 179 -203 188
rect -242 168 -211 170
rect -213 158 -211 168
rect -205 158 -203 175
rect -197 165 -195 188
rect -183 172 -174 176
rect -155 169 -153 172
rect -147 169 -145 172
rect -197 158 -195 161
rect -62 170 -60 188
rect -54 179 -52 188
rect -91 168 -60 170
rect -213 150 -211 153
rect -205 150 -203 153
rect -197 150 -195 153
rect -155 150 -153 159
rect -155 135 -153 146
rect -147 143 -145 159
rect -62 158 -60 168
rect -54 158 -52 175
rect -46 165 -44 188
rect -32 172 -23 176
rect -4 169 -2 172
rect 4 169 6 172
rect -46 158 -44 161
rect 78 170 80 188
rect 86 179 88 188
rect 49 168 80 170
rect -62 150 -60 153
rect -54 150 -52 153
rect -46 150 -44 153
rect -4 150 -2 159
rect -147 135 -145 139
rect -4 135 -2 146
rect 4 143 6 159
rect 78 158 80 168
rect 86 158 88 175
rect 94 165 96 188
rect 108 172 117 176
rect 136 169 138 172
rect 144 169 146 172
rect 94 158 96 161
rect 78 150 80 153
rect 86 150 88 153
rect 94 150 96 153
rect 136 150 138 159
rect 4 135 6 139
rect 136 135 138 146
rect 144 143 146 159
rect 161 143 163 153
rect 144 135 146 139
rect -155 127 -153 130
rect -147 127 -145 130
rect -4 127 -2 130
rect 4 127 6 130
rect 136 127 138 130
rect 144 127 146 130
rect -210 121 -208 124
rect -202 121 -200 124
rect -194 121 -192 124
rect -59 121 -57 124
rect -51 121 -49 124
rect -43 121 -41 124
rect 81 121 83 124
rect 89 121 91 124
rect 97 121 99 124
rect -210 84 -208 111
rect -202 98 -200 111
rect -202 84 -200 94
rect -194 91 -192 111
rect -157 104 -155 107
rect -149 104 -147 107
rect -141 104 -139 107
rect -194 84 -192 87
rect -157 85 -155 94
rect -210 76 -208 79
rect -202 76 -200 79
rect -194 75 -192 79
rect -157 64 -155 81
rect -149 78 -147 94
rect -149 64 -147 74
rect -141 71 -139 94
rect -59 84 -57 111
rect -51 98 -49 111
rect -51 84 -49 94
rect -43 91 -41 111
rect -6 104 -4 107
rect 2 104 4 107
rect 10 104 12 107
rect -43 84 -41 87
rect -6 85 -4 94
rect -59 76 -57 79
rect -51 76 -49 79
rect -43 75 -41 79
rect -141 64 -139 67
rect -6 64 -4 81
rect 2 78 4 94
rect 2 64 4 74
rect 10 71 12 94
rect 81 84 83 111
rect 89 98 91 111
rect 89 84 91 94
rect 97 91 99 111
rect 134 104 136 107
rect 142 104 144 107
rect 150 104 152 107
rect 97 84 99 87
rect 134 85 136 94
rect 81 76 83 79
rect 89 76 91 79
rect 97 75 99 79
rect 10 64 12 67
rect 134 64 136 81
rect 142 78 144 94
rect 142 64 144 74
rect 150 71 152 94
rect 150 64 152 67
rect -157 56 -155 59
rect -149 56 -147 59
rect -141 56 -139 59
rect -6 56 -4 59
rect 2 56 4 59
rect 10 56 12 59
rect 134 56 136 59
rect 142 56 144 59
rect 150 56 152 59
rect -212 53 -210 56
rect -204 53 -202 56
rect -196 53 -194 56
rect -61 53 -59 56
rect -53 53 -51 56
rect -45 53 -43 56
rect 79 53 81 56
rect 87 53 89 56
rect 95 53 97 56
rect -212 26 -210 43
rect -204 34 -202 43
rect -232 24 -210 26
rect -212 13 -210 24
rect -204 13 -202 30
rect -196 20 -194 43
rect -157 34 -155 37
rect -149 34 -147 37
rect -141 34 -139 37
rect -196 13 -194 16
rect -157 21 -155 24
rect -212 5 -210 8
rect -204 5 -202 8
rect -196 5 -194 8
rect -157 7 -155 17
rect -149 7 -147 24
rect -141 13 -139 24
rect -61 26 -59 43
rect -53 34 -51 43
rect -81 24 -59 26
rect -141 11 -104 13
rect -141 7 -139 11
rect -61 13 -59 24
rect -53 13 -51 30
rect -45 20 -43 43
rect 20 42 24 51
rect 3 28 5 31
rect 79 26 81 43
rect 87 34 89 43
rect 59 24 81 26
rect -45 13 -43 16
rect -61 5 -59 8
rect -53 5 -51 8
rect -45 5 -43 8
rect 3 6 5 18
rect 79 13 81 24
rect 87 13 89 30
rect 95 20 97 43
rect 160 42 164 51
rect 95 13 97 16
rect -157 -1 -155 2
rect -149 -9 -147 2
rect -141 -1 -139 2
rect 79 5 81 8
rect 87 5 89 8
rect 95 5 97 8
rect 3 -2 5 1
<< polycontact >>
rect -96 297 -92 301
rect -120 284 -116 288
rect 44 293 48 297
rect -82 287 -78 291
rect -96 268 -92 272
rect -232 247 -228 251
rect -212 240 -208 244
rect -232 233 -228 237
rect -204 233 -200 237
rect -145 248 -141 252
rect -153 227 -149 231
rect -137 241 -133 245
rect -129 234 -125 238
rect 59 287 63 291
rect 44 268 48 272
rect -61 240 -57 244
rect -81 233 -77 237
rect -53 233 -49 237
rect -1 230 3 234
rect 7 223 11 227
rect 79 240 83 244
rect 59 233 63 237
rect 87 233 91 237
rect 15 216 19 220
rect -246 167 -242 171
rect -207 175 -203 179
rect -187 172 -183 176
rect -174 172 -170 176
rect -199 161 -195 165
rect -95 167 -91 171
rect -56 175 -52 179
rect -157 146 -153 150
rect -36 172 -32 176
rect -23 172 -19 176
rect -48 161 -44 165
rect 45 167 49 171
rect 84 175 88 179
rect -6 146 -2 150
rect -149 139 -145 143
rect 104 172 108 176
rect 117 172 121 176
rect 92 161 96 165
rect 134 146 138 150
rect 2 139 6 143
rect 161 153 165 157
rect 142 139 146 143
rect 159 139 163 143
rect -214 101 -210 105
rect -204 94 -200 98
rect -63 101 -59 105
rect -196 87 -192 91
rect -159 81 -155 85
rect -151 74 -147 78
rect -53 94 -49 98
rect 77 101 81 105
rect -45 87 -41 91
rect -8 81 -4 85
rect -143 67 -139 71
rect 0 74 4 78
rect 87 94 91 98
rect 95 87 99 91
rect 132 81 136 85
rect 8 67 12 71
rect 140 74 144 78
rect 148 67 152 71
rect 20 51 24 55
rect -236 23 -232 27
rect -206 30 -202 34
rect -198 16 -194 20
rect -157 17 -153 21
rect -85 23 -81 27
rect -55 30 -51 34
rect -104 10 -100 14
rect 160 51 164 55
rect 20 38 24 42
rect -47 16 -43 20
rect 55 23 59 27
rect 85 30 89 34
rect -1 9 3 13
rect 160 38 164 42
rect 93 16 97 20
rect -150 -13 -146 -9
<< metal1 >>
rect -160 297 -96 300
rect -92 297 -72 300
rect -160 293 -157 297
rect -75 294 44 297
rect -227 290 -157 293
rect -154 291 -78 294
rect -227 257 -224 290
rect -154 287 -151 291
rect -245 254 -224 257
rect -221 284 -151 287
rect -78 287 59 290
rect -116 284 -99 287
rect -245 171 -242 254
rect -221 251 -218 284
rect -102 281 109 284
rect -162 278 -105 281
rect -211 268 -207 272
rect -203 268 -199 272
rect -215 263 -211 268
rect -199 263 -195 268
rect -235 247 -232 251
rect -228 248 -218 251
rect -207 250 -203 253
rect -162 252 -159 278
rect -108 275 103 278
rect -152 271 -148 275
rect -144 271 -140 275
rect -136 271 -132 275
rect -128 271 -124 275
rect -120 271 -116 275
rect -156 267 -152 271
rect -116 267 -112 271
rect -132 254 -128 257
rect -207 247 -194 250
rect -162 248 -145 252
rect -132 251 -119 254
rect -197 244 -194 247
rect -249 167 -246 171
rect -246 34 -242 167
rect -238 240 -212 244
rect -197 240 -177 244
rect -238 67 -235 240
rect -222 233 -204 237
rect -232 179 -229 233
rect -222 212 -218 233
rect -197 229 -194 240
rect -215 219 -211 224
rect -211 215 -207 219
rect -203 215 -199 219
rect -222 209 -183 212
rect -214 202 -210 206
rect -206 202 -202 206
rect -198 202 -194 206
rect -218 198 -214 202
rect -202 198 -198 202
rect -210 185 -206 188
rect -194 185 -190 188
rect -210 182 -190 185
rect -232 175 -207 179
rect -194 176 -190 182
rect -186 176 -183 209
rect -232 98 -229 175
rect -194 172 -187 176
rect -194 170 -189 172
rect -224 161 -199 165
rect -224 142 -221 161
rect -192 158 -189 170
rect -218 149 -214 153
rect -214 145 -210 149
rect -206 145 -202 149
rect -198 145 -194 149
rect -180 142 -177 240
rect -174 241 -137 245
rect -123 241 -119 251
rect -174 184 -171 241
rect -168 234 -129 238
rect -168 190 -165 234
rect -162 227 -153 231
rect -162 196 -159 227
rect -122 224 -119 241
rect -148 220 -128 223
rect -148 217 -144 220
rect -132 217 -128 220
rect -123 220 -106 224
rect -123 217 -119 220
rect -156 203 -152 212
rect -140 203 -136 212
rect -132 209 -128 212
rect -116 209 -112 212
rect -132 206 -112 209
rect -152 199 -148 203
rect -144 199 -140 203
rect -136 199 -132 203
rect -128 199 -124 203
rect -120 199 -116 203
rect -162 193 -121 196
rect -168 187 -127 190
rect -174 181 -133 184
rect -224 139 -177 142
rect -156 174 -152 178
rect -148 174 -144 178
rect -174 150 -171 172
rect -160 169 -156 174
rect -144 169 -140 174
rect -152 156 -148 159
rect -136 156 -133 181
rect -130 162 -127 187
rect -124 168 -121 193
rect -109 174 -106 220
rect -109 171 -98 174
rect -124 165 -104 168
rect -130 159 -110 162
rect -152 153 -139 156
rect -136 153 -116 156
rect -142 150 -139 153
rect -174 146 -157 150
rect -142 146 -122 150
rect -174 136 -171 146
rect -226 133 -171 136
rect -167 139 -149 143
rect -226 105 -223 133
rect -211 126 -207 130
rect -203 126 -199 130
rect -195 126 -191 130
rect -215 121 -211 126
rect -199 121 -195 126
rect -167 118 -163 139
rect -142 135 -139 146
rect -160 125 -156 130
rect -156 121 -152 125
rect -148 121 -144 125
rect -167 115 -128 118
rect -207 108 -203 111
rect -191 108 -187 111
rect -158 108 -154 112
rect -150 108 -146 112
rect -142 108 -138 112
rect -207 105 -186 108
rect -226 101 -214 105
rect -189 99 -186 105
rect -162 104 -158 108
rect -146 104 -142 108
rect -232 94 -204 98
rect -189 95 -177 99
rect -222 87 -196 91
rect -222 67 -218 87
rect -189 84 -186 95
rect -180 85 -177 95
rect -154 91 -150 94
rect -138 91 -134 94
rect -154 88 -134 91
rect -180 81 -159 85
rect -138 82 -134 88
rect -131 82 -128 115
rect -215 74 -211 79
rect -211 70 -207 74
rect -203 70 -199 74
rect -195 70 -191 74
rect -238 64 -183 67
rect -213 57 -209 61
rect -205 57 -201 61
rect -197 57 -193 61
rect -217 53 -213 57
rect -201 53 -197 57
rect -209 40 -205 43
rect -193 40 -189 43
rect -209 37 -189 40
rect -246 30 -206 34
rect -193 31 -189 37
rect -186 31 -183 64
rect -236 -15 -233 23
rect -229 -9 -226 30
rect -193 27 -183 31
rect -193 25 -188 27
rect -223 16 -198 20
rect -223 -3 -220 16
rect -191 13 -188 25
rect -217 4 -213 8
rect -213 0 -209 4
rect -205 0 -201 4
rect -197 0 -193 4
rect -180 -3 -177 81
rect -138 78 -128 82
rect -223 -6 -177 -3
rect -174 74 -151 78
rect -138 76 -133 78
rect -174 -9 -171 74
rect -168 67 -143 71
rect -168 48 -165 67
rect -136 64 -133 76
rect -162 55 -158 59
rect -158 51 -154 55
rect -150 51 -146 55
rect -142 51 -138 55
rect -125 48 -122 146
rect -168 45 -122 48
rect -158 38 -154 42
rect -150 38 -146 42
rect -142 38 -138 42
rect -138 34 -134 38
rect -165 13 -162 27
rect -119 21 -116 153
rect -153 17 -116 21
rect -165 10 -142 13
rect -229 -12 -171 -9
rect -168 7 -158 10
rect -146 7 -142 10
rect -168 -15 -165 7
rect -154 -2 -150 2
rect -138 -2 -134 2
rect -158 -6 -154 -2
rect -150 -6 -146 -2
rect -142 -6 -138 -2
rect -236 -18 -165 -15
rect -150 -33 -147 -13
rect -119 -27 -116 17
rect -113 -21 -110 159
rect -107 -15 -104 165
rect -101 27 -98 171
rect -95 171 -92 268
rect -60 268 -56 272
rect -52 268 -48 272
rect -64 263 -60 268
rect -48 263 -44 268
rect -56 250 -52 253
rect -56 247 -43 250
rect -46 244 -43 247
rect -87 240 -61 244
rect -46 240 -26 244
rect -95 34 -91 167
rect -87 67 -84 240
rect -71 233 -53 237
rect -81 179 -78 233
rect -71 212 -67 233
rect -46 229 -43 240
rect -64 219 -60 224
rect -60 215 -56 219
rect -52 215 -48 219
rect -71 209 -32 212
rect -63 202 -59 206
rect -55 202 -51 206
rect -47 202 -43 206
rect -67 198 -63 202
rect -51 198 -47 202
rect -59 185 -55 188
rect -43 185 -39 188
rect -59 182 -39 185
rect -81 175 -56 179
rect -43 176 -39 182
rect -35 176 -32 209
rect -81 98 -78 175
rect -43 172 -36 176
rect -43 170 -38 172
rect -73 161 -48 165
rect -73 142 -70 161
rect -41 158 -38 170
rect -67 149 -63 153
rect -63 145 -59 149
rect -55 145 -51 149
rect -47 145 -43 149
rect -29 142 -26 240
rect -10 234 -7 275
rect 0 259 4 263
rect 8 259 12 263
rect 16 259 20 263
rect 4 255 8 259
rect -4 241 0 245
rect 12 241 16 245
rect -4 238 16 241
rect 20 243 24 245
rect 20 237 25 243
rect -10 230 -1 234
rect -16 223 7 227
rect -16 184 -13 223
rect -10 216 15 220
rect -10 190 -7 216
rect 22 213 25 237
rect 12 212 25 213
rect 12 209 30 212
rect 12 206 16 209
rect -4 197 0 201
rect 20 197 24 201
rect 0 193 4 197
rect 8 193 12 197
rect 16 193 20 197
rect -10 187 24 190
rect -16 181 18 184
rect -73 139 -26 142
rect -5 174 -1 178
rect 3 174 7 178
rect -23 150 -20 172
rect -9 169 -5 174
rect 7 169 11 174
rect -1 156 3 159
rect -1 153 12 156
rect 9 150 12 153
rect 15 150 18 181
rect 21 156 24 187
rect 27 162 30 209
rect 45 171 48 268
rect 80 268 84 272
rect 88 268 92 272
rect 76 263 80 268
rect 92 263 96 268
rect 84 250 88 253
rect 100 250 103 275
rect 106 256 109 281
rect 106 253 126 256
rect 84 247 97 250
rect 100 247 120 250
rect 94 244 97 247
rect 53 240 79 244
rect 94 240 114 244
rect 27 159 42 162
rect 21 153 36 156
rect -23 146 -6 150
rect 9 146 30 150
rect -23 136 -20 146
rect -75 133 -20 136
rect -16 139 2 143
rect -75 105 -72 133
rect -60 126 -56 130
rect -52 126 -48 130
rect -44 126 -40 130
rect -64 121 -60 126
rect -48 121 -44 126
rect -16 118 -12 139
rect 9 135 12 146
rect -9 125 -5 130
rect -5 121 -1 125
rect 3 121 7 125
rect -16 115 23 118
rect -56 108 -52 111
rect -40 108 -36 111
rect -7 108 -3 112
rect 1 108 5 112
rect 9 108 13 112
rect -56 105 -35 108
rect -75 101 -63 105
rect -38 99 -35 105
rect -11 104 -7 108
rect 5 104 9 108
rect -81 94 -53 98
rect -38 95 -26 99
rect -71 87 -45 91
rect -71 67 -67 87
rect -38 84 -35 95
rect -29 85 -26 95
rect -3 91 1 94
rect 13 91 17 94
rect -3 88 17 91
rect -29 81 -8 85
rect 13 82 17 88
rect 20 82 23 115
rect 13 81 23 82
rect -64 74 -60 79
rect -60 70 -56 74
rect -52 70 -48 74
rect -44 70 -40 74
rect -87 64 -32 67
rect -62 57 -58 61
rect -54 57 -50 61
rect -46 57 -42 61
rect -66 53 -62 57
rect -50 53 -46 57
rect -58 40 -54 43
rect -42 40 -38 43
rect -58 37 -38 40
rect -95 30 -55 34
rect -42 31 -38 37
rect -35 31 -32 64
rect -101 24 -85 27
rect -78 -9 -75 30
rect -42 27 -32 31
rect -42 25 -37 27
rect -72 16 -47 20
rect -72 -3 -69 16
rect -40 13 -37 25
rect -66 4 -62 8
rect -62 0 -58 4
rect -54 0 -50 4
rect -46 0 -42 4
rect -29 -3 -26 81
rect 13 78 24 81
rect -72 -6 -26 -3
rect -23 74 0 78
rect 13 76 18 78
rect -23 -9 -20 74
rect -17 67 8 71
rect -17 48 -14 67
rect 15 64 18 76
rect -11 55 -7 59
rect 21 55 24 78
rect -7 51 -3 55
rect 1 51 5 55
rect 9 51 13 55
rect 27 48 30 146
rect -17 45 30 48
rect -78 -12 -20 -9
rect -17 39 20 42
rect -17 -15 -14 39
rect 2 32 6 36
rect 33 35 36 153
rect 16 32 36 35
rect -2 28 2 32
rect -107 -18 -14 -15
rect -11 9 -1 13
rect 6 12 10 18
rect 16 12 19 32
rect 39 27 42 159
rect 45 34 49 167
rect 53 67 56 240
rect 69 233 87 237
rect 59 179 62 233
rect 69 212 73 233
rect 94 229 97 240
rect 76 219 80 224
rect 80 215 84 219
rect 88 215 92 219
rect 69 209 108 212
rect 77 202 81 206
rect 85 202 89 206
rect 93 202 97 206
rect 73 198 77 202
rect 89 198 93 202
rect 81 185 85 188
rect 97 185 101 188
rect 81 182 101 185
rect 59 175 84 179
rect 97 176 101 182
rect 105 176 108 209
rect 59 98 62 175
rect 97 172 104 176
rect 97 170 102 172
rect 67 161 92 165
rect 67 142 70 161
rect 99 158 102 170
rect 73 149 77 153
rect 77 145 81 149
rect 85 145 89 149
rect 93 145 97 149
rect 111 142 114 240
rect 117 184 120 247
rect 123 190 126 253
rect 123 187 164 190
rect 117 181 158 184
rect 67 139 114 142
rect 135 174 139 178
rect 143 174 147 178
rect 117 150 120 172
rect 131 169 135 174
rect 147 169 151 174
rect 139 156 143 159
rect 139 153 152 156
rect 149 150 152 153
rect 155 150 158 181
rect 161 157 164 187
rect 117 146 134 150
rect 149 146 170 150
rect 117 136 120 146
rect 65 133 120 136
rect 124 139 142 143
rect 65 105 68 133
rect 80 126 84 130
rect 88 126 92 130
rect 96 126 100 130
rect 76 121 80 126
rect 92 121 96 126
rect 124 118 128 139
rect 149 135 152 146
rect 131 125 135 130
rect 135 121 139 125
rect 143 121 147 125
rect 160 118 163 139
rect 124 115 163 118
rect 84 108 88 111
rect 100 108 104 111
rect 133 108 137 112
rect 141 108 145 112
rect 149 108 153 112
rect 84 105 105 108
rect 65 101 77 105
rect 102 99 105 105
rect 129 104 133 108
rect 145 104 149 108
rect 59 94 87 98
rect 102 95 114 99
rect 69 87 95 91
rect 69 67 73 87
rect 102 84 105 95
rect 111 85 114 95
rect 137 91 141 94
rect 153 91 157 94
rect 137 88 157 91
rect 111 81 132 85
rect 153 82 157 88
rect 160 82 163 115
rect 153 81 163 82
rect 76 74 80 79
rect 80 70 84 74
rect 88 70 92 74
rect 96 70 100 74
rect 53 64 108 67
rect 78 57 82 61
rect 86 57 90 61
rect 94 57 98 61
rect 74 53 78 57
rect 90 53 94 57
rect 82 40 86 43
rect 98 40 102 43
rect 82 37 102 40
rect 45 30 85 34
rect 98 31 102 37
rect 105 31 108 64
rect 39 24 55 27
rect 6 9 19 12
rect -11 -21 -8 9
rect 6 6 10 9
rect -2 -3 2 1
rect 2 -7 6 -3
rect 13 -10 16 9
rect -113 -24 -8 -21
rect -5 -13 16 -10
rect 62 -9 65 30
rect 98 27 108 31
rect 98 25 103 27
rect 68 16 93 20
rect 68 -3 71 16
rect 100 13 103 25
rect 74 4 78 8
rect 78 0 82 4
rect 86 0 90 4
rect 94 0 98 4
rect 111 -3 114 81
rect 153 78 164 81
rect 68 -6 114 -3
rect 117 74 140 78
rect 153 76 158 78
rect 117 -9 120 74
rect 123 67 148 71
rect 123 48 126 67
rect 155 64 158 76
rect 129 55 133 59
rect 161 55 164 78
rect 133 51 137 55
rect 141 51 145 55
rect 149 51 153 55
rect 167 48 170 146
rect 123 45 170 48
rect 62 -12 120 -9
rect 123 39 160 42
rect -5 -27 -2 -13
rect 123 -15 126 39
rect 19 -16 126 -15
rect -119 -30 -2 -27
rect 1 -18 126 -16
rect 1 -19 22 -18
rect 1 -33 4 -19
rect -150 -36 4 -33
<< labels >>
rlabel nsubstratencontact -36 126 -36 130 1 Vdd!
rlabel psubstratepcontact -36 70 -36 74 1 GND!
rlabel psubstratepcontact 11 121 11 125 1 GND!
rlabel nsubstratencontact 11 174 11 178 1 Vdd!
rlabel nsubstratencontact -44 268 -44 272 1 Vdd!
rlabel psubstratepcontact -44 215 -44 219 1 GND!
rlabel nsubstratencontact -39 202 -39 206 1 Vdd!
rlabel psubstratepcontact -39 145 -39 149 1 GND!
rlabel nsubstratencontact -38 57 -38 61 1 Vdd!
rlabel psubstratepcontact -38 0 -38 4 1 GND!
rlabel nsubstratencontact 17 108 17 112 1 Vdd!
rlabel psubstratepcontact 17 51 17 55 1 GND!
rlabel metal1 23 80 23 85 1 QBNOT
rlabel metal1 30 76 30 84 1 QB
rlabel psubstratepcontact 10 -7 10 -3 1 GND!
rlabel nsubstratencontact 10 32 10 36 1 Vdd!
rlabel metal1 -10 9 -10 13 1 X
rlabel metal1 19 9 19 13 1 XNOT
rlabel nsubstratencontact -187 126 -187 130 1 Vdd!
rlabel psubstratepcontact -187 70 -187 74 1 GND!
rlabel psubstratepcontact -140 121 -140 125 1 GND!
rlabel nsubstratencontact -140 174 -140 178 1 Vdd!
rlabel nsubstratencontact -195 268 -195 272 1 Vdd!
rlabel psubstratepcontact -195 215 -195 219 1 GND!
rlabel nsubstratencontact -190 202 -190 206 1 Vdd!
rlabel psubstratepcontact -190 145 -190 149 1 GND!
rlabel nsubstratencontact -189 57 -189 61 1 Vdd!
rlabel psubstratepcontact -189 0 -189 4 1 GND!
rlabel nsubstratencontact -134 108 -134 112 1 Vdd!
rlabel psubstratepcontact -134 51 -134 55 1 GND!
rlabel metal1 -128 78 -128 83 1 QANOT
rlabel metal1 -122 78 -122 83 1 QA
rlabel nsubstratencontact -112 271 -112 275 1 Vdd!
rlabel nsubstratencontact -112 199 -112 203 1 GND!
rlabel nsubstratencontact -134 38 -134 42 1 Vdd!
rlabel psubstratepcontact -134 -6 -134 -2 1 GND!
rlabel nsubstratencontact 24 259 24 263 1 Vdd!
rlabel psubstratepcontact 24 193 24 197 1 GND!
rlabel nsubstratencontact 104 126 104 130 1 Vdd!
rlabel psubstratepcontact 104 70 104 74 1 GND!
rlabel psubstratepcontact 151 121 151 125 1 GND!
rlabel nsubstratencontact 151 174 151 178 1 Vdd!
rlabel nsubstratencontact 96 268 96 272 1 Vdd!
rlabel psubstratepcontact 96 215 96 219 1 GND!
rlabel nsubstratencontact 101 202 101 206 1 Vdd!
rlabel psubstratepcontact 101 145 101 149 1 GND!
rlabel nsubstratencontact 102 57 102 61 1 Vdd!
rlabel psubstratepcontact 102 0 102 4 1 GND!
rlabel nsubstratencontact 157 108 157 112 1 Vdd!
rlabel psubstratepcontact 157 51 157 55 1 GND!
rlabel metal1 163 78 163 85 1 QCNOT
rlabel metal1 170 78 170 85 1 QC
rlabel metal1 -235 247 -235 251 1 CLK
rlabel metal1 -249 167 -249 171 3 RESET
rlabel polycontact -236 23 -236 27 1 inA
rlabel polycontact -85 23 -85 27 1 inB
rlabel polycontact 55 23 55 27 1 inC
rlabel space -160 -14 -160 -10 1 gateForAflipFlop
rlabel space -113 234 -113 239 1 gateForBflipFlop
rlabel space 28 222 29 228 1 gateForCflipFlop
rlabel metal1 -119 17 -119 21 1 xNotForA
rlabel polycontact -146 -13 -146 -9 1 cNotForA
rlabel polycontact -100 10 -100 14 1 bNotForA
rlabel metal1 -10 230 -10 234 1 cForC
rlabel metal1 -16 223 -16 227 1 bForC
rlabel metal1 -10 216 -10 220 1 xNotForC
rlabel metal1 25 209 25 212 1 cGateOut
rlabel metal1 -168 7 -168 10 1 aGateOut
rlabel metal1 -106 219 -106 224 1 bGateOut
rlabel metal1 -162 248 -162 252 1 cForB
rlabel metal1 -174 240 -174 245 1 xNotForB
rlabel metal1 -168 233 -168 238 1 xForB
rlabel metal1 -162 226 -162 231 1 bNotForB
rlabel polycontact -120 284 -120 288 1 cNotForB
<< end >>
