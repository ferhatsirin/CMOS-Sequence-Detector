magic
tech scmos
timestamp 1578763967
<< nwell >>
rect 46 113 79 142
rect 43 47 83 75
rect 101 19 134 48
rect 46 -29 86 0
rect 99 -47 139 -19
rect 44 -98 84 -70
<< polysilicon >>
rect 57 129 59 132
rect 65 129 67 132
rect 57 110 59 119
rect 57 95 59 106
rect 65 103 67 119
rect 65 95 67 99
rect 57 87 59 90
rect 65 87 67 90
rect 54 64 56 67
rect 62 64 64 67
rect 70 64 72 67
rect 26 41 35 45
rect 54 36 56 54
rect 62 45 64 54
rect 25 34 56 36
rect 54 24 56 34
rect 62 24 64 41
rect 70 31 72 54
rect 84 38 93 42
rect 112 35 114 38
rect 120 35 122 38
rect 70 24 72 27
rect 54 16 56 19
rect 62 16 64 19
rect 70 16 72 19
rect 112 16 114 25
rect 112 1 114 12
rect 120 9 122 25
rect 120 1 122 5
rect 112 -7 114 -4
rect 120 -7 122 -4
rect 57 -13 59 -10
rect 65 -13 67 -10
rect 73 -13 75 -10
rect 57 -50 59 -23
rect 65 -36 67 -23
rect 65 -50 67 -40
rect 73 -43 75 -23
rect 110 -30 112 -27
rect 118 -30 120 -27
rect 126 -30 128 -27
rect 73 -50 75 -47
rect 110 -49 112 -40
rect 57 -58 59 -55
rect 65 -58 67 -55
rect 73 -59 75 -55
rect 110 -70 112 -53
rect 118 -56 120 -40
rect 118 -70 120 -60
rect 126 -63 128 -40
rect 139 -56 148 -52
rect 126 -70 128 -67
rect 110 -78 112 -75
rect 118 -78 120 -75
rect 126 -78 128 -75
rect 55 -81 57 -78
rect 63 -81 65 -78
rect 71 -81 73 -78
rect 55 -108 57 -91
rect 63 -100 65 -91
rect 35 -110 57 -108
rect 55 -121 57 -110
rect 63 -121 65 -104
rect 71 -114 73 -91
rect 71 -121 73 -118
rect 55 -129 57 -126
rect 63 -129 65 -126
rect 71 -129 73 -126
<< ndiffusion >>
rect 56 90 57 95
rect 59 90 65 95
rect 67 90 68 95
rect 53 19 54 24
rect 56 19 62 24
rect 64 19 70 24
rect 72 19 73 24
rect 111 -4 112 1
rect 114 -4 120 1
rect 122 -4 123 1
rect 56 -55 57 -50
rect 59 -55 65 -50
rect 67 -55 73 -50
rect 75 -55 76 -50
rect 109 -75 110 -70
rect 112 -75 118 -70
rect 120 -75 126 -70
rect 128 -75 129 -70
rect 54 -126 55 -121
rect 57 -126 63 -121
rect 65 -126 71 -121
rect 73 -126 74 -121
<< pdiffusion >>
rect 56 119 57 129
rect 59 119 60 129
rect 64 119 65 129
rect 67 119 68 129
rect 53 54 54 64
rect 56 54 57 64
rect 61 54 62 64
rect 64 54 65 64
rect 69 54 70 64
rect 72 54 73 64
rect 111 25 112 35
rect 114 25 115 35
rect 119 25 120 35
rect 122 25 123 35
rect 56 -23 57 -13
rect 59 -23 60 -13
rect 64 -23 65 -13
rect 67 -23 68 -13
rect 72 -23 73 -13
rect 75 -23 76 -13
rect 109 -40 110 -30
rect 112 -40 113 -30
rect 117 -40 118 -30
rect 120 -40 121 -30
rect 125 -40 126 -30
rect 128 -40 129 -30
rect 54 -91 55 -81
rect 57 -91 58 -81
rect 62 -91 63 -81
rect 65 -91 66 -81
rect 70 -91 71 -81
rect 73 -91 74 -81
<< metal1 >>
rect 56 134 60 138
rect 64 134 68 138
rect 52 129 56 134
rect 68 129 72 134
rect 60 116 64 119
rect 60 113 73 116
rect 70 110 73 113
rect 29 106 55 110
rect 70 106 90 110
rect 21 -100 25 33
rect 29 -67 32 106
rect 45 99 63 103
rect 45 78 49 99
rect 70 95 73 106
rect 52 85 56 90
rect 56 81 60 85
rect 64 81 68 85
rect 45 75 84 78
rect 53 68 57 72
rect 61 68 65 72
rect 69 68 73 72
rect 49 64 53 68
rect 65 64 69 68
rect 57 51 61 54
rect 73 51 77 54
rect 57 48 77 51
rect 39 41 60 45
rect 73 42 77 48
rect 81 42 84 75
rect 35 -36 38 41
rect 73 38 80 42
rect 73 36 78 38
rect 43 27 68 31
rect 43 8 46 27
rect 75 24 78 36
rect 49 15 53 19
rect 53 11 57 15
rect 61 11 65 15
rect 69 11 73 15
rect 87 8 90 106
rect 43 5 90 8
rect 111 40 115 44
rect 119 40 123 44
rect 93 16 96 38
rect 107 35 111 40
rect 123 35 127 40
rect 115 22 119 25
rect 115 19 128 22
rect 125 16 128 19
rect 93 12 110 16
rect 125 12 145 16
rect 93 2 96 12
rect 41 -1 96 2
rect 100 5 118 9
rect 41 -29 44 -1
rect 56 -8 60 -4
rect 64 -8 68 -4
rect 72 -8 76 -4
rect 52 -13 56 -8
rect 68 -13 72 -8
rect 100 -16 104 5
rect 125 1 128 12
rect 107 -9 111 -4
rect 111 -13 115 -9
rect 119 -13 123 -9
rect 100 -19 139 -16
rect 60 -26 64 -23
rect 76 -26 80 -23
rect 109 -26 113 -22
rect 117 -26 121 -22
rect 125 -26 129 -22
rect 60 -29 81 -26
rect 41 -33 53 -29
rect 78 -35 81 -29
rect 105 -30 109 -26
rect 121 -30 125 -26
rect 35 -40 63 -36
rect 78 -39 90 -35
rect 45 -47 71 -43
rect 45 -67 49 -47
rect 78 -50 81 -39
rect 87 -49 90 -39
rect 113 -43 117 -40
rect 129 -43 133 -40
rect 113 -46 133 -43
rect 87 -53 108 -49
rect 129 -52 133 -46
rect 136 -52 139 -19
rect 52 -60 56 -55
rect 56 -64 60 -60
rect 64 -64 68 -60
rect 72 -64 76 -60
rect 29 -70 84 -67
rect 54 -77 58 -73
rect 62 -77 66 -73
rect 70 -77 74 -73
rect 50 -81 54 -77
rect 66 -81 70 -77
rect 58 -94 62 -91
rect 74 -94 78 -91
rect 58 -97 78 -94
rect 21 -104 61 -100
rect 74 -103 78 -97
rect 81 -103 84 -70
rect 29 -111 31 -107
rect 38 -143 41 -104
rect 74 -107 84 -103
rect 74 -109 79 -107
rect 44 -118 69 -114
rect 44 -137 47 -118
rect 76 -121 79 -109
rect 50 -130 54 -126
rect 54 -134 58 -130
rect 62 -134 66 -130
rect 70 -134 74 -130
rect 87 -137 90 -53
rect 129 -56 135 -52
rect 142 -38 145 12
rect 142 -42 151 -38
rect 44 -140 90 -137
rect 93 -60 116 -56
rect 129 -58 134 -56
rect 93 -143 96 -60
rect 99 -67 124 -63
rect 99 -86 102 -67
rect 131 -70 134 -58
rect 105 -79 109 -75
rect 109 -83 113 -79
rect 117 -83 121 -79
rect 125 -83 129 -79
rect 142 -86 145 -42
rect 152 -56 156 -52
rect 99 -89 145 -86
rect 38 -146 96 -143
<< ntransistor >>
rect 57 90 59 95
rect 65 90 67 95
rect 54 19 56 24
rect 62 19 64 24
rect 70 19 72 24
rect 112 -4 114 1
rect 120 -4 122 1
rect 57 -55 59 -50
rect 65 -55 67 -50
rect 73 -55 75 -50
rect 110 -75 112 -70
rect 118 -75 120 -70
rect 126 -75 128 -70
rect 55 -126 57 -121
rect 63 -126 65 -121
rect 71 -126 73 -121
<< ptransistor >>
rect 57 119 59 129
rect 65 119 67 129
rect 54 54 56 64
rect 62 54 64 64
rect 70 54 72 64
rect 112 25 114 35
rect 120 25 122 35
rect 57 -23 59 -13
rect 65 -23 67 -13
rect 73 -23 75 -13
rect 110 -40 112 -30
rect 118 -40 120 -30
rect 126 -40 128 -30
rect 55 -91 57 -81
rect 63 -91 65 -81
rect 71 -91 73 -81
<< polycontact >>
rect 55 106 59 110
rect 63 99 67 103
rect 22 41 26 45
rect 35 41 39 45
rect 21 33 25 37
rect 60 41 64 45
rect 80 38 84 42
rect 93 38 97 42
rect 68 27 72 31
rect 110 12 114 16
rect 118 5 122 9
rect 53 -33 57 -29
rect 63 -40 67 -36
rect 71 -47 75 -43
rect 108 -53 112 -49
rect 116 -60 120 -56
rect 135 -56 139 -52
rect 148 -56 152 -52
rect 124 -67 128 -63
rect 31 -111 35 -107
rect 61 -104 65 -100
rect 69 -118 73 -114
<< ndcontact >>
rect 52 90 56 95
rect 68 90 73 95
rect 49 19 53 24
rect 73 19 78 24
rect 107 -4 111 1
rect 123 -4 128 1
rect 52 -55 56 -50
rect 76 -55 81 -50
rect 105 -75 109 -70
rect 129 -75 134 -70
rect 50 -126 54 -121
rect 74 -126 79 -121
<< pdcontact >>
rect 52 119 56 129
rect 60 119 64 129
rect 68 119 72 129
rect 49 54 53 64
rect 57 54 61 64
rect 65 54 69 64
rect 73 54 77 64
rect 107 25 111 35
rect 115 25 119 35
rect 123 25 127 35
rect 52 -23 56 -13
rect 60 -23 64 -13
rect 68 -23 72 -13
rect 76 -23 80 -13
rect 105 -40 109 -30
rect 113 -40 117 -30
rect 121 -40 125 -30
rect 129 -40 133 -30
rect 50 -91 54 -81
rect 58 -91 62 -81
rect 66 -91 70 -81
rect 74 -91 78 -81
<< psubstratepcontact >>
rect 52 81 56 85
rect 60 81 64 85
rect 68 81 72 85
rect 49 11 53 15
rect 57 11 61 15
rect 65 11 69 15
rect 73 11 77 15
rect 107 -13 111 -9
rect 115 -13 119 -9
rect 123 -13 127 -9
rect 52 -64 56 -60
rect 60 -64 64 -60
rect 68 -64 72 -60
rect 76 -64 80 -60
rect 105 -83 109 -79
rect 113 -83 117 -79
rect 121 -83 125 -79
rect 129 -83 133 -79
rect 50 -134 54 -130
rect 58 -134 62 -130
rect 66 -134 70 -130
rect 74 -134 78 -130
<< nsubstratencontact >>
rect 52 134 56 138
rect 60 134 64 138
rect 68 134 72 138
rect 49 68 53 72
rect 57 68 61 72
rect 65 68 69 72
rect 73 68 77 72
rect 107 40 111 44
rect 115 40 119 44
rect 123 40 127 44
rect 52 -8 56 -4
rect 60 -8 64 -4
rect 68 -8 72 -4
rect 76 -8 80 -4
rect 105 -26 109 -22
rect 113 -26 117 -22
rect 121 -26 125 -22
rect 129 -26 133 -22
rect 50 -77 54 -73
rect 58 -77 62 -73
rect 66 -77 70 -73
rect 74 -77 78 -73
<< labels >>
rlabel nsubstratencontact 80 -8 80 -4 1 Vdd!
rlabel psubstratepcontact 80 -64 80 -60 1 GND!
rlabel psubstratepcontact 127 -13 127 -9 1 GND!
rlabel nsubstratencontact 127 40 127 44 1 Vdd!
rlabel nsubstratencontact 72 134 72 138 1 Vdd!
rlabel psubstratepcontact 72 81 72 85 1 GND!
rlabel nsubstratencontact 77 68 77 72 1 Vdd!
rlabel psubstratepcontact 77 11 77 15 1 GND!
rlabel polycontact 22 41 22 45 3 CLK
rlabel polycontact 21 33 21 37 3 RESET
rlabel nsubstratencontact 78 -77 78 -73 1 Vdd!
rlabel psubstratepcontact 78 -134 78 -130 1 GND!
rlabel nsubstratencontact 133 -26 133 -22 1 Vdd!
rlabel psubstratepcontact 133 -83 133 -79 1 GND!
rlabel metal1 156 -56 156 -52 7 QNOT
rlabel metal1 151 -42 151 -38 7 Q
rlabel metal1 29 -111 29 -107 1 D
<< end >>
