magic
tech scmos
timestamp 1578774135
<< nwell >>
rect 73 57 113 84
<< polysilicon >>
rect 84 73 86 76
rect 92 73 94 76
rect 100 73 102 76
rect 84 60 86 63
rect 84 46 86 56
rect 92 46 94 63
rect 100 46 102 63
rect 84 38 86 41
rect 92 30 94 41
rect 100 38 102 41
<< ndiffusion >>
rect 83 41 84 46
rect 86 41 87 46
rect 91 41 92 46
rect 94 41 95 46
rect 99 41 100 46
rect 102 41 103 46
<< pdiffusion >>
rect 83 63 84 73
rect 86 63 92 73
rect 94 63 100 73
rect 102 63 103 73
<< metal1 >>
rect 83 77 87 81
rect 91 77 95 81
rect 99 77 103 81
rect 103 73 107 77
rect 76 52 79 66
rect 88 56 115 60
rect 76 49 99 52
rect 73 46 83 49
rect 95 46 99 49
rect 87 37 91 41
rect 103 37 107 41
rect 83 33 87 37
rect 91 33 95 37
rect 99 33 103 37
<< ntransistor >>
rect 84 41 86 46
rect 92 41 94 46
rect 100 41 102 46
<< ptransistor >>
rect 84 63 86 73
rect 92 63 94 73
rect 100 63 102 73
<< polycontact >>
rect 84 56 88 60
rect 102 49 106 53
rect 91 26 95 30
<< ndcontact >>
rect 79 41 83 46
rect 87 41 91 46
rect 95 41 99 46
rect 103 41 107 46
<< pdcontact >>
rect 79 63 83 73
rect 103 63 107 73
<< psubstratepcontact >>
rect 79 33 83 37
rect 87 33 91 37
rect 95 33 99 37
rect 103 33 107 37
<< nsubstratencontact >>
rect 79 77 83 81
rect 87 77 91 81
rect 95 77 99 81
rect 103 77 107 81
<< labels >>
rlabel nsubstratencontact 107 77 107 81 1 Vdd!
rlabel psubstratepcontact 107 33 107 37 1 GND!
rlabel polycontact 95 26 95 30 1 cNotForA
rlabel metal1 73 46 73 49 1 aGateOut
rlabel metal1 115 56 115 60 1 xNotForA
rlabel polycontact 106 49 106 53 1 bNotForA
<< end >>
