magic
tech scmos
timestamp 1578831393
<< nwell >>
rect 78 291 135 318
<< ntransistor >>
rect 89 252 91 257
rect 97 252 99 257
rect 105 252 107 257
rect 113 252 115 257
rect 121 252 123 257
<< ptransistor >>
rect 89 297 91 307
rect 97 297 99 307
rect 105 297 107 307
rect 113 297 115 307
rect 121 297 123 307
<< ndiffusion >>
rect 88 252 89 257
rect 91 252 92 257
rect 96 252 97 257
rect 99 252 100 257
rect 104 252 105 257
rect 107 252 108 257
rect 112 252 113 257
rect 115 252 116 257
rect 120 252 121 257
rect 123 252 124 257
<< pdiffusion >>
rect 88 297 89 307
rect 91 297 97 307
rect 99 297 105 307
rect 107 297 108 307
rect 112 297 113 307
rect 115 297 121 307
rect 123 297 124 307
<< ndcontact >>
rect 84 252 88 257
rect 92 252 96 257
rect 100 252 104 257
rect 108 252 112 257
rect 116 252 120 257
rect 124 252 128 257
<< pdcontact >>
rect 84 297 88 307
rect 108 297 112 307
rect 124 297 128 307
<< nsubstratencontact >>
rect 84 311 88 315
rect 92 311 96 315
rect 100 311 104 315
rect 108 311 112 315
rect 116 311 120 315
rect 124 311 128 315
rect 84 239 88 243
rect 92 239 96 243
rect 100 239 104 243
rect 108 239 112 243
rect 116 239 120 243
rect 124 239 128 243
<< polysilicon >>
rect 89 307 91 310
rect 97 307 99 310
rect 105 307 107 310
rect 113 307 115 310
rect 121 307 123 320
rect 89 271 91 297
rect 97 292 99 297
rect 89 257 91 267
rect 97 257 99 288
rect 105 285 107 297
rect 105 257 107 281
rect 113 278 115 297
rect 113 257 115 274
rect 121 257 123 297
rect 89 249 91 252
rect 97 249 99 252
rect 105 249 107 252
rect 113 249 115 252
rect 121 249 123 252
<< polycontact >>
rect 120 320 124 324
rect 95 288 99 292
rect 87 267 91 271
rect 103 281 107 285
rect 111 274 115 278
<< metal1 >>
rect 88 311 92 315
rect 96 311 100 315
rect 104 311 108 315
rect 112 311 116 315
rect 120 311 124 315
rect 84 307 88 311
rect 124 307 128 311
rect 108 294 112 297
rect 78 288 95 292
rect 108 291 121 294
rect 66 281 103 285
rect 117 281 121 291
rect 72 274 111 278
rect 78 267 87 271
rect 118 264 121 281
rect 92 260 112 263
rect 92 257 96 260
rect 108 257 112 260
rect 117 260 134 264
rect 117 257 121 260
rect 84 243 88 252
rect 100 243 104 252
rect 108 249 112 252
rect 124 249 128 252
rect 108 246 128 249
rect 88 239 92 243
rect 96 239 100 243
rect 104 239 108 243
rect 112 239 116 243
rect 120 239 124 243
<< labels >>
rlabel nsubstratencontact 128 311 128 315 1 Vdd!
rlabel nsubstratencontact 128 239 128 243 1 GND!
rlabel metal1 78 288 78 292 1 cForB
rlabel polycontact 120 320 120 324 1 cNotForB
rlabel metal1 66 281 66 285 3 xNotForB
rlabel metal1 72 274 72 278 1 xForB
rlabel metal1 78 267 78 271 1 bNotForB
rlabel metal1 134 260 134 264 7 bGateOut
<< end >>
