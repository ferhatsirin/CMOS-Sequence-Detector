magic
tech scmos
timestamp 1578774809
<< nwell >>
rect 228 278 270 305
<< ntransistor >>
rect 240 240 242 245
rect 248 240 250 245
rect 256 240 258 245
<< ptransistor >>
rect 240 284 242 294
rect 248 284 250 294
rect 256 284 258 294
<< ndiffusion >>
rect 239 240 240 245
rect 242 240 248 245
rect 250 240 251 245
rect 255 240 256 245
rect 258 240 259 245
<< pdiffusion >>
rect 239 284 240 294
rect 242 284 243 294
rect 247 284 248 294
rect 250 284 251 294
rect 255 284 256 294
rect 258 284 259 294
<< ndcontact >>
rect 235 240 239 245
rect 251 240 255 245
rect 259 240 263 245
<< pdcontact >>
rect 235 284 239 294
rect 243 284 247 294
rect 251 284 255 294
rect 259 284 263 294
<< psubstratepcontact >>
rect 235 232 239 236
rect 243 232 247 236
rect 251 232 255 236
rect 259 232 263 236
<< nsubstratencontact >>
rect 235 298 239 302
rect 243 298 247 302
rect 251 298 255 302
rect 259 298 263 302
<< polysilicon >>
rect 240 294 242 297
rect 248 294 250 297
rect 256 294 258 297
rect 240 273 242 284
rect 240 245 242 269
rect 248 266 250 284
rect 248 245 250 262
rect 256 259 258 284
rect 256 245 258 255
rect 240 237 242 240
rect 248 237 250 240
rect 256 237 258 240
<< polycontact >>
rect 238 269 242 273
rect 246 262 250 266
rect 254 255 258 259
<< metal1 >>
rect 239 298 243 302
rect 247 298 251 302
rect 255 298 259 302
rect 243 294 247 298
rect 235 280 239 284
rect 251 280 255 284
rect 235 277 255 280
rect 259 282 263 284
rect 259 276 264 282
rect 229 269 238 273
rect 223 262 246 266
rect 229 255 254 259
rect 261 252 264 276
rect 251 248 264 252
rect 251 245 255 248
rect 235 236 239 240
rect 259 236 263 240
rect 239 232 243 236
rect 247 232 251 236
rect 255 232 259 236
<< labels >>
rlabel nsubstratencontact 263 298 263 302 1 Vdd!
rlabel psubstratepcontact 263 232 263 236 1 GND!
rlabel metal1 229 269 229 273 1 cForC
rlabel metal1 223 262 223 266 1 bForC
rlabel metal1 229 255 229 259 1 xNotForC
rlabel metal1 264 248 264 251 1 cGateOut
<< end >>
